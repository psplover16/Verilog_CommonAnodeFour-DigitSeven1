module tt(clk,seg,way,showDigit,showNum);
input clk;// 
output reg[7:0] seg;
output reg[7:0] way; 
// 
input [3:0] showDigit; 
input [5:0] showNum;
// 
reg[21:0] frequency;
// reg [5:0] tmpshowNum;
// 
reg[5:0] aaa;
// assign way = showDigit; // 秀第幾位數
// 
always@(posedge clk)frequency=frequency+1;   
// 


always @(posedge showDigit or posedge showNum or posedge showNum[5])begin

    case(showDigit)

       1: way = 8'b00000001;
       2: way = 8'b00000010;
       3: way = 8'b00000100;
       4: way = 8'b00001000;
       5: way = 8'b00010000;
       6: way = 8'b00100000;
       7: way = 8'b01000000;
       8: way = 8'b10000000;
       default: way = 8'b11111111; // 8.
    endcase


    case(showNum)

      0: seg = 8'b01111110;
      1: seg = 8'b00110000;
      2: seg = 8'b01101101;
      3: seg = 8'b01111001;
      4: seg = 8'b00110011;
      5: seg = 8'b01011011;
      6: seg = 8'b01011111;
      7: seg = 8'b01110010;
      8: seg = 8'b01111111;
      9: seg = 8'b11110011;
      default: seg = 8'b11111111; // 8.
    endcase

// 
if(showNum[5]==1)seg[0] = 1;


end
endmodule

